
library IEEE;
use IEEE.STD_Logic_1164.all;

entity BCD is
	port(
	bcd_in: in std_Logic_Vector(3 downto 0);
	seven_seg: out std_Logic_Vector(6 downto 0)
	);
end BCD;

architecture comportamento of BCD is
begin
	
	 with bcd_in select 
        seven_seg <= "1000000" when "0000",
             "1111001" when "0001", 
             "0100100" when "0010",       
             "0110000" when "0011",       
             "0011001" when "0100",       
             "0010010" when "0101",       
             "0000010" when "0110",       
             "1111000" when "0111",       
             "0000000" when "1000",       
             "0010000" when "1001",       
             "0001000" when "1010",       
             "0000011" when "1011",       
             "1000110" when "1100",       
             "0100001" when "1101",       
             "0000110" when "1110",       
             "0001110" when others; 
	
end comportamento;